* I:\3. East West University\BSC   IN   CSE\COURSE\5th SEMESTER = SUMMER 2021\CSE209\CSE209 Lab Experiment\Lab 6\class task.sch

* Schematics Version 9.1 - Web Update 1
* Mon Sep 06 15:28:03 2021


.PARAM         RVAR=10 

** Analysis setup **
.DC LIN PARAM RVAR 1 2000 0.1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "class task.net"
.INC "class task.als"


.probe


.END
