* I:\3. East West University\BSC   IN   CSE\COURSE\5th SEMESTER = SUMMER 2021\CSE209\CSE209 Lab Experiment\Project\Project.sch

* Schematics Version 9.1 - Web Update 1
* Wed Sep 08 15:21:36 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Project.net"
.INC "Project.als"


.probe


.END
