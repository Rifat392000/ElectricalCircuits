* I:\3. East West University\BSC   IN   CSE\COURSE\5th SEMESTER = SUMMER 2021\CSE209\CSE209 Lab Experiment\Lab 6\Lab Material\Experiment 6.sch

* Schematics Version 9.1 - Web Update 1
* Sat Sep 11 16:45:48 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Experiment 6.net"
.INC "Experiment 6.als"


.probe


.END
