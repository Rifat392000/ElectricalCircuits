* I:\3. East West University\BSC   IN   CSE\COURSE\5th SEMESTER = SUMMER 2021\CSE209\CSE209 Lab Experiment\Lab 7\Experiment 7 part1.sch

* Schematics Version 9.1 - Web Update 1
* Mon Sep 06 09:40:23 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Experiment 7 part1.net"
.INC "Experiment 7 part1.als"


.probe


.END
