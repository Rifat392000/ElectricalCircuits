* I:\3. East West University\BSC   IN   CSE\COURSE\5th SEMESTER = SUMMER 2021\CSE209\CSE209 Lab Experiment\Lab 7\Experiment 7 part4.sch

* Schematics Version 9.1 - Web Update 1
* Wed Sep 08 16:33:01 2021


.PARAM         RVAR=10 

** Analysis setup **
.DC LIN PARAM RVAR 1 20 0.1 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Experiment 7 part4.net"
.INC "Experiment 7 part4.als"


.probe


.END
