* I:\3. East West University\BSC   IN   CSE\COURSE\5th SEMESTER = SUMMER 2021\CSE209\CSE209 Lab Experiment\Lab 7\Experiment 7 part2.sch

* Schematics Version 9.1 - Web Update 1
* Mon Sep 06 09:53:57 2021



** Analysis setup **
.DC LIN V_E 0V 20V 1V 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Experiment 7 part2.net"
.INC "Experiment 7 part2.als"


.probe


.END
